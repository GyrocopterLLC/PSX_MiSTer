module cpu_top
(
    input  clk1x,
    input  clk2x,
    input  clk3x,
    input  ce,
    input  reset,
    input  TURBO,
    input  TURBO_CACHE,
    input  TURBO_CACHE50,
    input  irqRequest,
    input  dmaStallCPU,
    input  cpuPaused,
    output error,
    output error2,
    output mem_request,
    output mem_rnw,
    output mem_isData,
    output mem_isCache,
    output [3:0] mem_oldtagvalids,
    output [31:0] mem_addressInstr,
    output [31:0] mem_addressData,
    output [1:0] mem_reqsize,
    output [3:0] mem_writeMask,
    output [31:0] mem_dataWrite,
    input  [31:0] mem_dataRead,
    input  mem_done,
    input  mem_fifofull,
    input  [3:0] mem_tagvalids,
    input  [3:0] cache_wr,
    input  [31:0] cache_data,
    input  [7:0] cache_addr,
    output stallNext,
    input  [20:0] dma_cache_Adr,
    input  [31:0] dma_cache_data,
    input  dma_cache_write,
    input  ram_done,
    input  ram_rnw,
    input  [31:0] ram_dataRead,
    input  gte_busy,
    output gte_readEna,
    output [5:0] gte_readAddr,
    input  [31:0] gte_readData,
    output [5:0] gte_writeAddr,
    output [31:0] gte_writeData,
    output gte_writeEna,
    output [31:0] gte_cmdData,
    output gte_cmdEna,
    input  SS_reset,
    input  [31:0] SS_DataWrite,
    input  [7:0] SS_Adr,
    input  SS_wren_CPU,
    input  SS_wren_SCP,
    input  SS_rden_CPU,
    input  SS_rden_SCP,
    output [31:0] SS_DataRead_CPU,
    output [31:0] SS_DataRead_SCP,
    output SS_idle,
    input  debug_firstGTE
    
);

sdram_model3x my_sdram(
    .clk(clk1x),
    .clk3x,
    .refresh(reset_intern),
    .addr({2'b00, ram_Adr}),
    .req(ram_ena),
    .ram_dma(ram_dma),
    .ram_dmacnt(ram_cntDMA),
    .ram_iscache(ram_iscache),
    .rnw(ram_rnw),
    .be(ram_be),
    .di(ram_dataWrite),
    .dout(),
    .do32(ram_dataRead32),
    .done(ram_done),
    .cache_wr(cache_wr),
    .cache_data(cache_data),
    .cache_addr(cache_addr),
    .dma_wr(dma_wr),
    .dma_data(dma_data),
    .reqprocessed(dma_reqprocessed),
    .ram_idle(),
    .ram_dmafifo_adr(ram_dmafifo_adr),
    .ram_dmafifo_data (ram_dmafifo_data),
    .ram_dmafifo_empty(ram_dmafifo_empty),
    .ram_dmafifo_read(ram_dmafifo_read)
);

cpu my_cpu(
    .clk1x,
    .clk2x,
    .clk3x,
    .ce,
    .reset,
    .TURBO,
    .TURBO_CACHE,
    .TURBO_CACHE50,
    .irqRequest,
    .dmaStallCPU,
    .cpuPaused,
    .error,
    .error2,
    .mem_request,
    .mem_rnw,
    .mem_isData,
    .mem_isCache,
    .mem_oldtagvalids,
    .mem_addressInstr,
    .mem_addressData,
    .mem_reqsize,
    .mem_writeMask,
    .mem_dataWrite,
    .mem_dataRead,
    .mem_done,
    .mem_fifofull,
    .mem_tagvalids,
    .cache_wr,
    .cache_data,
    .cache_addr,
    .stallNext,
    .dma_cache_Adr,
    .dma_cache_data,
    .dma_cache_write,
    .ram_done,
    .ram_rnw,
    .ram_dataRead,
    .gte_busy,
    .gte_readEna,
    .gte_readAddr,
    .gte_readData,
    .gte_writeAddr,
    .gte_writeData,
    .gte_writeEna,
    .gte_cmdData,
    .gte_cmdEna,
    .SS_reset,
    .SS_DataWrite,
    .SS_Adr,
    .SS_wren_CPU,
    .SS_wren_SCP,
    .SS_rden_CPU,
    .SS_rden_SCP,
    .SS_DataRead_CPU,
    .SS_DataRead_SCP,
    .SS_idle,
    .debug_firstGTE
);

endmodule

